module chip_7458 ( // Описание модуля, реализующего логику И-НЕ 7458
    p1a, p1b, p1c, p1d, p1e, p1f, // Входы первой группы (две тройки для двух 3-входовых И)
    p1y, // Выход первой группы (ИЛИ из двух 3-входовых И)
    p2a, p2b, p2c, p2d, // Входы второй группы (две пары для двух 2-входовых И)
    p2y ); // Выход второй группы (ИЛИ из двух 2-входовых И)

input p1a, p1b, p1c, p1d, p1e, p1f; // Объявление входов первой группы
input p2a, p2b, p2c, p2d; // Объявление входов второй группы
output p1y; // Объявление выхода первой группы
output p2y; // Объявление выхода второй группы

assign p1y = (p1a & p1b & p1c) | (p1d & p1e & p1f); // Первая функция: (A&B&C) OR (D&E&F)
assign p2y = (p2a & p2b) | (p2c & p2d); // Вторая функция: (A&B) OR (C&D)

endmodule // Конец описания модуля